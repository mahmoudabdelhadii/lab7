`define MNONE 2'b00 //do not read or write
`define MWRITE 2'b01 // write to memory(can change)
`define MREAD  2'b11 // read from memory(can change)
module MEM(/*INPUTS*/clk,mem_cmd,mem_addr,write_data, /*OUTPUTS*/read_data );
input clk;
input[15:0] write_data;
output[15:0] read_data;
input [1:0] mem_cmd;
input [8:0] mem_addr;

wire [15:0] tribufferin;

wire msel;
wire[15:0] mwriteeq,mreadeq;
wire writeout,readout;
assign msel = (mem_addr[8:8] == 1'b0)? 1'b1: 1'b0;
RAM #(16,8) MEMORY(.clk(clk),.read_address(mem_addr[7:0]),.write_address(mem_addr[7:0]),.write(writeout),.din(write_data),.dout(tribufferin));


assign mwriteeq = (mem_cmd == `MWRITE)? 1'b1: 1'b0;
assign mreadeq  = (mem_cmd == `MREAD)? 1'b1: 1'b0;

assign writeout = mwriteeq & msel;
assign readout = mreadeq &msel;

tristate_buffer#(16) tribuf(tribufferin, readout, read_data);


endmodule
module RAM(clk,read_address,write_address,write,din,dout);
  parameter data_width = 32; 
  parameter addr_width = 4;
  parameter filename = "data.txt";

  input clk;
  input [addr_width-1:0] read_address, write_address;
  input write;
  input [data_width-1:0] din;
  output [data_width-1:0] dout;
  reg [data_width-1:0] dout;

  reg [data_width-1:0] mem [2**addr_width-1:0];

  initial $readmemb(filename, mem);

  always @ (posedge clk) begin
    if (write)
      mem[write_address] <= din;
    dout <= mem[read_address]; // dout doesn't get din in this clock cycle 
                               // (this is due to Verilog non-blocking assignment "<=")
  end 
endmodule