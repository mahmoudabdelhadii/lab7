module PC(/*inputs*/load_pc, reset_pc, load_addr, addr_sel,datapath_out,/*outputs*/read_data,write_data,mem_addr,mem_cmd);
input


